module lightpwm_tb();

endmodule
