module light-pwm(
  // system
  input clk,

  // sensor
  output sensor_ncs,
  output sensor_scl,
  input  sensor_sda,
  
  // rgb-led
  output led0_r,
  output led0_g,
  output led0_b,
);

endmodule

