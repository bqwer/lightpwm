module filter(
  input        clk,
  input  [7:0] sensor_data,
  output [7:0] mean_data
};

endmodule

