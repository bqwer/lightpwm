module color (
  input  [7:0] sensor_data,

  output [7:0] red_pwm,
  output [7:0] green_pwm,
  output [7:0] blue_pwm,
);

endmodule

