module (
  input        clk,
  output       sensor_ncs,
  output       sensor_scl,
  input        sensor_sda
  output [7:0] sensor_data,
)

endmodule
